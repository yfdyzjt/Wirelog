module Input_Single (       
    input wire in,
    output wire out
);
    
    assign out = in;

endmodule