module Output_Single_Wire (       
    input wire in,
    output wire out
);
    
    assign out = in;

endmodule